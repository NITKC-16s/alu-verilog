module NOT1 (
	input A,
	output X );

    assign X = ~A;

endmodule


module NOT1 (
	input A,
	output X );

	NAND2 new_nand (A,A, X);

endmodule
